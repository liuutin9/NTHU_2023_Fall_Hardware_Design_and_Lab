`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/10/06 08:47:11
// Design Name: 
// Module Name: Lab2_111060013_Carry_Look_Ahead_Adder_8bit_t
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Lab2_111060013_Carry_Look_Ahead_Adder_8bit_t(

    );
endmodule
